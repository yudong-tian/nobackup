netcdf lis_input.clm45 {
dimensions:
        east_west = 288 ;
        north_south = 192 ;
        east_west_b = 292 ;
        north_south_b = 196 ;
        east_west_GDAS_T126 = 384 ;
        north_south_GDAS_T126 = 190 ;
        east_west_GDAS_T170 = 512 ;
        north_south_GDAS_T170 = 256 ;
        east_west_GDAS_T254 = 768 ;
        north_south_GDAS_T254 = 384 ;
        east_west_GDAS_T382 = 1152 ;
        north_south_GDAS_T382 = 576 ;
        east_west_GDAS_T574 = 1760 ;
        north_south_GDAS_T574 = 880 ;
        east_west_GDAS_T1534 = 3072 ;
        north_south_GDAS_T1534 = 1536 ;
        month = 12 ;
        time = 1 ;
        sfctypes = 14 ;
        soilfracbins = 1 ;
        elevbins = 1 ;

        ncorners = 4; 

	nglcec = 10 ;
	nglcecp1 = 11 ;
	numurbl = 3 ;
	nlevurb = 5 ;
	numrad = 2 ;
	nchar = 256 ;
	nlevsoi = 10 ;
	lsmpft = 17 ;

variables:
        float time(time) ;
  double xc(north_south, east_west) ;
                xc:standard_name = "xc" ;
                xc:units = "" ;
                xc:scale_factor = 1.f ;
                xc:add_offset = 0.f ;
                xc:missing_value = -9999.f ;
                xc:vmin = 0.f ;
                xc:vmax = 0.f ;
                xc:num_bins = 1 ;
  double yc(north_south, east_west) ;
                yc:standard_name = "yc" ;
                yc:units = "" ;
                yc:scale_factor = 1.f ;
                yc:add_offset = 0.f ;
                yc:missing_value = -9999.f ;
                yc:vmin = 0.f ;
                yc:vmax = 0.f ;
                yc:num_bins = 1 ;
  double xv(north_south, east_west, ncorners) ;
                xv:standard_name = "xv" ;
                xv:units = "" ;
                xv:scale_factor = 1.f ;
                xv:add_offset = 0.f ;
                xv:missing_value = -9999.f ;
                xv:vmin = 0.f ;
                xv:vmax = 0.f ;
                xv:num_bins = 1 ;
  double yv(north_south, east_west, ncorners) ;
                yv:standard_name = "yv" ;
                yv:units = "" ;
                yv:scale_factor = 1.f ;
                yv:add_offset = 0.f ;
                yv:missing_value = -9999.f ;
                yv:vmin = 0.f ;
                yv:vmax = 0.f ;
                yv:num_bins = 1 ;
  int LANDMASK(north_south, east_west) ;
                LANDMASK:standard_name = "LANDMASK" ;
                LANDMASK:units = "" ;
                LANDMASK:scale_factor = 1.f ;
                LANDMASK:add_offset = 0.f ;
                LANDMASK:missing_value = -9999.f ;
                LANDMASK:vmin = 0.f ;
                LANDMASK:vmax = 0.f ;
                LANDMASK:num_bins = 1 ;
  double area(north_south, east_west) ;
                area:standard_name = "area" ;
                area:units = "" ;
                area:scale_factor = 1.f ;
                area:add_offset = 0.f ;
                area:missing_value = -9999.f ;
                area:vmin = 0.f ;
                area:vmax = 0.f ;
                area:num_bins = 1 ;
  double frac(north_south, east_west) ;
                frac:standard_name = "frac" ;
                frac:units = "" ;
                frac:scale_factor = 1.f ;
                frac:add_offset = 0.f ;
                frac:missing_value = -9999.f ;
                frac:vmin = 0.f ;
                frac:vmax = 0.f ;
                frac:num_bins = 1 ;
  int mxsoil_color ;
                mxsoil_color:standard_name = "mxsoil_color" ;
                mxsoil_color:units = "" ;
                mxsoil_color:scale_factor = 1.f ;
                mxsoil_color:add_offset = 0.f ;
                mxsoil_color:missing_value = -9999.f ;
                mxsoil_color:vmin = 0.f ;
                mxsoil_color:vmax = 0.f ;
                mxsoil_color:num_bins = 1 ;
  int SOIL_COLOR(north_south, east_west) ;
                SOIL_COLOR:standard_name = "SOIL_COLOR" ;
                SOIL_COLOR:units = "" ;
                SOIL_COLOR:scale_factor = 1.f ;
                SOIL_COLOR:add_offset = 0.f ;
                SOIL_COLOR:missing_value = -9999.f ;
                SOIL_COLOR:vmin = 0.f ;
                SOIL_COLOR:vmax = 0.f ;
                SOIL_COLOR:num_bins = 1 ;
  double PCT_SAND(nlevsoi, north_south, east_west) ;
                PCT_SAND:standard_name = "PCT_SAND" ;
                PCT_SAND:units = "" ;
                PCT_SAND:scale_factor = 1.f ;
                PCT_SAND:add_offset = 0.f ;
                PCT_SAND:missing_value = -9999.f ;
                PCT_SAND:vmin = 0.f ;
                PCT_SAND:vmax = 0.f ;
                PCT_SAND:num_bins = 1 ;
  double PCT_CLAY(nlevsoi, north_south, east_west) ;
                PCT_CLAY:standard_name = "PCT_CLAY" ;
                PCT_CLAY:units = "" ;
                PCT_CLAY:scale_factor = 1.f ;
                PCT_CLAY:add_offset = 0.f ;
                PCT_CLAY:missing_value = -9999.f ;
                PCT_CLAY:vmin = 0.f ;
                PCT_CLAY:vmax = 0.f ;
                PCT_CLAY:num_bins = 1 ;
  double ORGANIC(nlevsoi, north_south, east_west) ;
                ORGANIC:standard_name = "ORGANIC" ;
                ORGANIC:units = "" ;
                ORGANIC:scale_factor = 1.f ;
                ORGANIC:add_offset = 0.f ;
                ORGANIC:missing_value = -9999.f ;
                ORGANIC:vmin = 0.f ;
                ORGANIC:vmax = 0.f ;
                ORGANIC:num_bins = 1 ;
  double FMAX(north_south, east_west) ;
                FMAX:standard_name = "FMAX" ;
                FMAX:units = "" ;
                FMAX:scale_factor = 1.f ;
                FMAX:add_offset = 0.f ;
                FMAX:missing_value = -9999.f ;
                FMAX:vmin = 0.f ;
                FMAX:vmax = 0.f ;
                FMAX:num_bins = 1 ;
  double LANDFRAC_PFT(north_south, east_west) ;
                LANDFRAC_PFT:standard_name = "LANDFRAC_PFT" ;
                LANDFRAC_PFT:units = "" ;
                LANDFRAC_PFT:scale_factor = 1.f ;
                LANDFRAC_PFT:add_offset = 0.f ;
                LANDFRAC_PFT:missing_value = -9999.f ;
                LANDFRAC_PFT:vmin = 0.f ;
                LANDFRAC_PFT:vmax = 0.f ;
                LANDFRAC_PFT:num_bins = 1 ;
  int PFTDATA_MASK(north_south, east_west) ;
                PFTDATA_MASK:standard_name = "PFTDATA_MASK" ;
                PFTDATA_MASK:units = "" ;
                PFTDATA_MASK:scale_factor = 1.f ;
                PFTDATA_MASK:add_offset = 0.f ;
                PFTDATA_MASK:missing_value = -9999.f ;
                PFTDATA_MASK:vmin = 0.f ;
                PFTDATA_MASK:vmax = 0.f ;
                PFTDATA_MASK:num_bins = 1 ;
  double PCT_PFT(lsmpft, north_south, east_west) ;
                PCT_PFT:standard_name = "PCT_PFT" ;
                PCT_PFT:units = "" ;
                PCT_PFT:scale_factor = 1.f ;
                PCT_PFT:add_offset = 0.f ;
                PCT_PFT:missing_value = -9999.f ;
                PCT_PFT:vmin = 0.f ;
                PCT_PFT:vmax = 0.f ;
                PCT_PFT:num_bins = 1 ;
  double MONTHLY_LAI(month, lsmpft, north_south, east_west) ;
                MONTHLY_LAI:standard_name = "MONTHLY_LAI" ;
                MONTHLY_LAI:units = "" ;
                MONTHLY_LAI:scale_factor = 1.f ;
                MONTHLY_LAI:add_offset = 0.f ;
                MONTHLY_LAI:missing_value = -9999.f ;
                MONTHLY_LAI:vmin = 0.f ;
                MONTHLY_LAI:vmax = 0.f ;
                MONTHLY_LAI:num_bins = 1 ;
  double MONTHLY_SAI(month, lsmpft, north_south, east_west) ;
                MONTHLY_SAI:standard_name = "MONTHLY_SAI" ;
                MONTHLY_SAI:units = "" ;
                MONTHLY_SAI:scale_factor = 1.f ;
                MONTHLY_SAI:add_offset = 0.f ;
                MONTHLY_SAI:missing_value = -9999.f ;
                MONTHLY_SAI:vmin = 0.f ;
                MONTHLY_SAI:vmax = 0.f ;
                MONTHLY_SAI:num_bins = 1 ;
  double MONTHLY_HEIGHT_TOP(month, lsmpft, north_south, east_west) ;
                MONTHLY_HEIGHT_TOP:standard_name = "MONTHLY_HEIGHT_TOP" ;
                MONTHLY_HEIGHT_TOP:units = "" ;
                MONTHLY_HEIGHT_TOP:scale_factor = 1.f ;
                MONTHLY_HEIGHT_TOP:add_offset = 0.f ;
                MONTHLY_HEIGHT_TOP:missing_value = -9999.f ;
                MONTHLY_HEIGHT_TOP:vmin = 0.f ;
                MONTHLY_HEIGHT_TOP:vmax = 0.f ;
                MONTHLY_HEIGHT_TOP:num_bins = 1 ;
  double MONTHLY_HEIGHT_BOT(month, lsmpft, north_south, east_west) ;
                MONTHLY_HEIGHT_BOT:standard_name = "MONTHLY_HEIGHT_BOT" ;
                MONTHLY_HEIGHT_BOT:units = "" ;
                MONTHLY_HEIGHT_BOT:scale_factor = 1.f ;
                MONTHLY_HEIGHT_BOT:add_offset = 0.f ;
                MONTHLY_HEIGHT_BOT:missing_value = -9999.f ;
                MONTHLY_HEIGHT_BOT:vmin = 0.f ;
                MONTHLY_HEIGHT_BOT:vmax = 0.f ;
                MONTHLY_HEIGHT_BOT:num_bins = 1 ;
  int month(month) ;
                month:standard_name = "month" ;
                month:units = "" ;
                month:scale_factor = 1.f ;
                month:add_offset = 0.f ;
                month:missing_value = -9999.f ;
                month:vmin = 0.f ;
                month:vmax = 0.f ;
                month:num_bins = 1 ;
  double AREA(north_south, east_west) ;
                AREA:standard_name = "AREA" ;
                AREA:units = "" ;
                AREA:scale_factor = 1.f ;
                AREA:add_offset = 0.f ;
                AREA:missing_value = -9999.f ;
                AREA:vmin = 0.f ;
                AREA:vmax = 0.f ;
                AREA:num_bins = 1 ;
  double LONGXY(north_south, east_west) ;
                LONGXY:standard_name = "LONGXY" ;
                LONGXY:units = "" ;
                LONGXY:scale_factor = 1.f ;
                LONGXY:add_offset = 0.f ;
                LONGXY:missing_value = -9999.f ;
                LONGXY:vmin = 0.f ;
                LONGXY:vmax = 0.f ;
                LONGXY:num_bins = 1 ;
  double LATIXY(north_south, east_west) ;
                LATIXY:standard_name = "LATIXY" ;
                LATIXY:units = "" ;
                LATIXY:scale_factor = 1.f ;
                LATIXY:add_offset = 0.f ;
                LATIXY:missing_value = -9999.f ;
                LATIXY:vmin = 0.f ;
                LATIXY:vmax = 0.f ;
                LATIXY:num_bins = 1 ;
  double EF1_BTR(north_south, east_west) ;
                EF1_BTR:standard_name = "EF1_BTR" ;
                EF1_BTR:units = "" ;
                EF1_BTR:scale_factor = 1.f ;
                EF1_BTR:add_offset = 0.f ;
                EF1_BTR:missing_value = -9999.f ;
                EF1_BTR:vmin = 0.f ;
                EF1_BTR:vmax = 0.f ;
                EF1_BTR:num_bins = 1 ;
  double EF1_FET(north_south, east_west) ;
                EF1_FET:standard_name = "EF1_FET" ;
                EF1_FET:units = "" ;
                EF1_FET:scale_factor = 1.f ;
                EF1_FET:add_offset = 0.f ;
                EF1_FET:missing_value = -9999.f ;
                EF1_FET:vmin = 0.f ;
                EF1_FET:vmax = 0.f ;
                EF1_FET:num_bins = 1 ;
  double EF1_FDT(north_south, east_west) ;
                EF1_FDT:standard_name = "EF1_FDT" ;
                EF1_FDT:units = "" ;
                EF1_FDT:scale_factor = 1.f ;
                EF1_FDT:add_offset = 0.f ;
                EF1_FDT:missing_value = -9999.f ;
                EF1_FDT:vmin = 0.f ;
                EF1_FDT:vmax = 0.f ;
                EF1_FDT:num_bins = 1 ;
  double EF1_SHR(north_south, east_west) ;
                EF1_SHR:standard_name = "EF1_SHR" ;
                EF1_SHR:units = "" ;
                EF1_SHR:scale_factor = 1.f ;
                EF1_SHR:add_offset = 0.f ;
                EF1_SHR:missing_value = -9999.f ;
                EF1_SHR:vmin = 0.f ;
                EF1_SHR:vmax = 0.f ;
                EF1_SHR:num_bins = 1 ;
  double EF1_GRS(north_south, east_west) ;
                EF1_GRS:standard_name = "EF1_GRS" ;
                EF1_GRS:units = "" ;
                EF1_GRS:scale_factor = 1.f ;
                EF1_GRS:add_offset = 0.f ;
                EF1_GRS:missing_value = -9999.f ;
                EF1_GRS:vmin = 0.f ;
                EF1_GRS:vmax = 0.f ;
                EF1_GRS:num_bins = 1 ;
  double EF1_CRP(north_south, east_west) ;
                EF1_CRP:standard_name = "EF1_CRP" ;
                EF1_CRP:units = "" ;
                EF1_CRP:scale_factor = 1.f ;
                EF1_CRP:add_offset = 0.f ;
                EF1_CRP:missing_value = -9999.f ;
                EF1_CRP:vmin = 0.f ;
                EF1_CRP:vmax = 0.f ;
                EF1_CRP:num_bins = 1 ;
  double CANYON_HWR(numurbl, north_south, east_west) ;
                CANYON_HWR:standard_name = "CANYON_HWR" ;
                CANYON_HWR:units = "" ;
                CANYON_HWR:scale_factor = 1.f ;
                CANYON_HWR:add_offset = 0.f ;
                CANYON_HWR:missing_value = -9999.f ;
                CANYON_HWR:vmin = 0.f ;
                CANYON_HWR:vmax = 0.f ;
                CANYON_HWR:num_bins = 1 ;
  double EM_IMPROAD(numurbl, north_south, east_west) ;
                EM_IMPROAD:standard_name = "EM_IMPROAD" ;
                EM_IMPROAD:units = "" ;
                EM_IMPROAD:scale_factor = 1.f ;
                EM_IMPROAD:add_offset = 0.f ;
                EM_IMPROAD:missing_value = -9999.f ;
                EM_IMPROAD:vmin = 0.f ;
                EM_IMPROAD:vmax = 0.f ;
                EM_IMPROAD:num_bins = 1 ;
  double EM_PERROAD(numurbl, north_south, east_west) ;
                EM_PERROAD:standard_name = "EM_PERROAD" ;
                EM_PERROAD:units = "" ;
                EM_PERROAD:scale_factor = 1.f ;
                EM_PERROAD:add_offset = 0.f ;
                EM_PERROAD:missing_value = -9999.f ;
                EM_PERROAD:vmin = 0.f ;
                EM_PERROAD:vmax = 0.f ;
                EM_PERROAD:num_bins = 1 ;
  double EM_ROOF(numurbl, north_south, east_west) ;
                EM_ROOF:standard_name = "EM_ROOF" ;
                EM_ROOF:units = "" ;
                EM_ROOF:scale_factor = 1.f ;
                EM_ROOF:add_offset = 0.f ;
                EM_ROOF:missing_value = -9999.f ;
                EM_ROOF:vmin = 0.f ;
                EM_ROOF:vmax = 0.f ;
                EM_ROOF:num_bins = 1 ;
  double EM_WALL(numurbl, north_south, east_west) ;
                EM_WALL:standard_name = "EM_WALL" ;
                EM_WALL:units = "" ;
                EM_WALL:scale_factor = 1.f ;
                EM_WALL:add_offset = 0.f ;
                EM_WALL:missing_value = -9999.f ;
                EM_WALL:vmin = 0.f ;
                EM_WALL:vmax = 0.f ;
                EM_WALL:num_bins = 1 ;
  double HT_ROOF(numurbl, north_south, east_west) ;
                HT_ROOF:standard_name = "HT_ROOF" ;
                HT_ROOF:units = "" ;
                HT_ROOF:scale_factor = 1.f ;
                HT_ROOF:add_offset = 0.f ;
                HT_ROOF:missing_value = -9999.f ;
                HT_ROOF:vmin = 0.f ;
                HT_ROOF:vmax = 0.f ;
                HT_ROOF:num_bins = 1 ;
  double THICK_ROOF(numurbl, north_south, east_west) ;
                THICK_ROOF:standard_name = "THICK_ROOF" ;
                THICK_ROOF:units = "" ;
                THICK_ROOF:scale_factor = 1.f ;
                THICK_ROOF:add_offset = 0.f ;
                THICK_ROOF:missing_value = -9999.f ;
                THICK_ROOF:vmin = 0.f ;
                THICK_ROOF:vmax = 0.f ;
                THICK_ROOF:num_bins = 1 ;
  double THICK_WALL(numurbl, north_south, east_west) ;
                THICK_WALL:standard_name = "THICK_WALL" ;
                THICK_WALL:units = "" ;
                THICK_WALL:scale_factor = 1.f ;
                THICK_WALL:add_offset = 0.f ;
                THICK_WALL:missing_value = -9999.f ;
                THICK_WALL:vmin = 0.f ;
                THICK_WALL:vmax = 0.f ;
                THICK_WALL:num_bins = 1 ;
  double T_BUILDING_MAX(numurbl, north_south, east_west) ;
                T_BUILDING_MAX:standard_name = "T_BUILDING_MAX" ;
                T_BUILDING_MAX:units = "" ;
                T_BUILDING_MAX:scale_factor = 1.f ;
                T_BUILDING_MAX:add_offset = 0.f ;
                T_BUILDING_MAX:missing_value = -9999.f ;
                T_BUILDING_MAX:vmin = 0.f ;
                T_BUILDING_MAX:vmax = 0.f ;
                T_BUILDING_MAX:num_bins = 1 ;
  double T_BUILDING_MIN(numurbl, north_south, east_west) ;
                T_BUILDING_MIN:standard_name = "T_BUILDING_MIN" ;
                T_BUILDING_MIN:units = "" ;
                T_BUILDING_MIN:scale_factor = 1.f ;
                T_BUILDING_MIN:add_offset = 0.f ;
                T_BUILDING_MIN:missing_value = -9999.f ;
                T_BUILDING_MIN:vmin = 0.f ;
                T_BUILDING_MIN:vmax = 0.f ;
                T_BUILDING_MIN:num_bins = 1 ;
  double WIND_HGT_CANYON(numurbl, north_south, east_west) ;
                WIND_HGT_CANYON:standard_name = "WIND_HGT_CANYON" ;
                WIND_HGT_CANYON:units = "" ;
                WIND_HGT_CANYON:scale_factor = 1.f ;
                WIND_HGT_CANYON:add_offset = 0.f ;
                WIND_HGT_CANYON:missing_value = -9999.f ;
                WIND_HGT_CANYON:vmin = 0.f ;
                WIND_HGT_CANYON:vmax = 0.f ;
                WIND_HGT_CANYON:num_bins = 1 ;
  double WTLUNIT_ROOF(numurbl, north_south, east_west) ;
                WTLUNIT_ROOF:standard_name = "WTLUNIT_ROOF" ;
                WTLUNIT_ROOF:units = "" ;
                WTLUNIT_ROOF:scale_factor = 1.f ;
                WTLUNIT_ROOF:add_offset = 0.f ;
                WTLUNIT_ROOF:missing_value = -9999.f ;
                WTLUNIT_ROOF:vmin = 0.f ;
                WTLUNIT_ROOF:vmax = 0.f ;
                WTLUNIT_ROOF:num_bins = 1 ;
  double WTROAD_PERV(numurbl, north_south, east_west) ;
                WTROAD_PERV:standard_name = "WTROAD_PERV" ;
                WTROAD_PERV:units = "" ;
                WTROAD_PERV:scale_factor = 1.f ;
                WTROAD_PERV:add_offset = 0.f ;
                WTROAD_PERV:missing_value = -9999.f ;
                WTROAD_PERV:vmin = 0.f ;
                WTROAD_PERV:vmax = 0.f ;
                WTROAD_PERV:num_bins = 1 ;
  double ALB_IMPROAD_DIR(numrad, numurbl, north_south, east_west) ;
                ALB_IMPROAD_DIR:standard_name = "ALB_IMPROAD_DIR" ;
                ALB_IMPROAD_DIR:units = "" ;
                ALB_IMPROAD_DIR:scale_factor = 1.f ;
                ALB_IMPROAD_DIR:add_offset = 0.f ;
                ALB_IMPROAD_DIR:missing_value = -9999.f ;
                ALB_IMPROAD_DIR:vmin = 0.f ;
                ALB_IMPROAD_DIR:vmax = 0.f ;
                ALB_IMPROAD_DIR:num_bins = 1 ;
  double ALB_IMPROAD_DIF(numrad, numurbl, north_south, east_west) ;
                ALB_IMPROAD_DIF:standard_name = "ALB_IMPROAD_DIF" ;
                ALB_IMPROAD_DIF:units = "" ;
                ALB_IMPROAD_DIF:scale_factor = 1.f ;
                ALB_IMPROAD_DIF:add_offset = 0.f ;
                ALB_IMPROAD_DIF:missing_value = -9999.f ;
                ALB_IMPROAD_DIF:vmin = 0.f ;
                ALB_IMPROAD_DIF:vmax = 0.f ;
                ALB_IMPROAD_DIF:num_bins = 1 ;
  double ALB_PERROAD_DIR(numrad, numurbl, north_south, east_west) ;
                ALB_PERROAD_DIR:standard_name = "ALB_PERROAD_DIR" ;
                ALB_PERROAD_DIR:units = "" ;
                ALB_PERROAD_DIR:scale_factor = 1.f ;
                ALB_PERROAD_DIR:add_offset = 0.f ;
                ALB_PERROAD_DIR:missing_value = -9999.f ;
                ALB_PERROAD_DIR:vmin = 0.f ;
                ALB_PERROAD_DIR:vmax = 0.f ;
                ALB_PERROAD_DIR:num_bins = 1 ;
  double ALB_PERROAD_DIF(numrad, numurbl, north_south, east_west) ;
                ALB_PERROAD_DIF:standard_name = "ALB_PERROAD_DIF" ;
                ALB_PERROAD_DIF:units = "" ;
                ALB_PERROAD_DIF:scale_factor = 1.f ;
                ALB_PERROAD_DIF:add_offset = 0.f ;
                ALB_PERROAD_DIF:missing_value = -9999.f ;
                ALB_PERROAD_DIF:vmin = 0.f ;
                ALB_PERROAD_DIF:vmax = 0.f ;
                ALB_PERROAD_DIF:num_bins = 1 ;
  double ALB_ROOF_DIR(numrad, numurbl, north_south, east_west) ;
                ALB_ROOF_DIR:standard_name = "ALB_ROOF_DIR" ;
                ALB_ROOF_DIR:units = "" ;
                ALB_ROOF_DIR:scale_factor = 1.f ;
                ALB_ROOF_DIR:add_offset = 0.f ;
                ALB_ROOF_DIR:missing_value = -9999.f ;
                ALB_ROOF_DIR:vmin = 0.f ;
                ALB_ROOF_DIR:vmax = 0.f ;
                ALB_ROOF_DIR:num_bins = 1 ;
  double ALB_ROOF_DIF(numrad, numurbl, north_south, east_west) ;
                ALB_ROOF_DIF:standard_name = "ALB_ROOF_DIF" ;
                ALB_ROOF_DIF:units = "" ;
                ALB_ROOF_DIF:scale_factor = 1.f ;
                ALB_ROOF_DIF:add_offset = 0.f ;
                ALB_ROOF_DIF:missing_value = -9999.f ;
                ALB_ROOF_DIF:vmin = 0.f ;
                ALB_ROOF_DIF:vmax = 0.f ;
                ALB_ROOF_DIF:num_bins = 1 ;
  double ALB_WALL_DIR(numrad, numurbl, north_south, east_west) ;
                ALB_WALL_DIR:standard_name = "ALB_WALL_DIR" ;
                ALB_WALL_DIR:units = "" ;
                ALB_WALL_DIR:scale_factor = 1.f ;
                ALB_WALL_DIR:add_offset = 0.f ;
                ALB_WALL_DIR:missing_value = -9999.f ;
                ALB_WALL_DIR:vmin = 0.f ;
                ALB_WALL_DIR:vmax = 0.f ;
                ALB_WALL_DIR:num_bins = 1 ;
  double ALB_WALL_DIF(numrad, numurbl, north_south, east_west) ;
                ALB_WALL_DIF:standard_name = "ALB_WALL_DIF" ;
                ALB_WALL_DIF:units = "" ;
                ALB_WALL_DIF:scale_factor = 1.f ;
                ALB_WALL_DIF:add_offset = 0.f ;
                ALB_WALL_DIF:missing_value = -9999.f ;
                ALB_WALL_DIF:vmin = 0.f ;
                ALB_WALL_DIF:vmax = 0.f ;
                ALB_WALL_DIF:num_bins = 1 ;
  double TK_ROOF(nlevurb, numurbl, north_south, east_west) ;
                TK_ROOF:standard_name = "TK_ROOF" ;
                TK_ROOF:units = "" ;
                TK_ROOF:scale_factor = 1.f ;
                TK_ROOF:add_offset = 0.f ;
                TK_ROOF:missing_value = -9999.f ;
                TK_ROOF:vmin = 0.f ;
                TK_ROOF:vmax = 0.f ;
                TK_ROOF:num_bins = 1 ;
  double TK_WALL(nlevurb, numurbl, north_south, east_west) ;
                TK_WALL:standard_name = "TK_WALL" ;
                TK_WALL:units = "" ;
                TK_WALL:scale_factor = 1.f ;
                TK_WALL:add_offset = 0.f ;
                TK_WALL:missing_value = -9999.f ;
                TK_WALL:vmin = 0.f ;
                TK_WALL:vmax = 0.f ;
                TK_WALL:num_bins = 1 ;
  double TK_IMPROAD(nlevurb, numurbl, north_south, east_west) ;
                TK_IMPROAD:standard_name = "TK_IMPROAD" ;
                TK_IMPROAD:units = "" ;
                TK_IMPROAD:scale_factor = 1.f ;
                TK_IMPROAD:add_offset = 0.f ;
                TK_IMPROAD:missing_value = -9999.f ;
                TK_IMPROAD:vmin = 0.f ;
                TK_IMPROAD:vmax = 0.f ;
                TK_IMPROAD:num_bins = 1 ;
  double CV_ROOF(nlevurb, numurbl, north_south, east_west) ;
                CV_ROOF:standard_name = "CV_ROOF" ;
                CV_ROOF:units = "" ;
                CV_ROOF:scale_factor = 1.f ;
                CV_ROOF:add_offset = 0.f ;
                CV_ROOF:missing_value = -9999.f ;
                CV_ROOF:vmin = 0.f ;
                CV_ROOF:vmax = 0.f ;
                CV_ROOF:num_bins = 1 ;
  double CV_WALL(nlevurb, numurbl, north_south, east_west) ;
                CV_WALL:standard_name = "CV_WALL" ;
                CV_WALL:units = "" ;
                CV_WALL:scale_factor = 1.f ;
                CV_WALL:add_offset = 0.f ;
                CV_WALL:missing_value = -9999.f ;
                CV_WALL:vmin = 0.f ;
                CV_WALL:vmax = 0.f ;
                CV_WALL:num_bins = 1 ;
  double CV_IMPROAD(nlevurb, numurbl, north_south, east_west) ;
                CV_IMPROAD:standard_name = "CV_IMPROAD" ;
                CV_IMPROAD:units = "" ;
                CV_IMPROAD:scale_factor = 1.f ;
                CV_IMPROAD:add_offset = 0.f ;
                CV_IMPROAD:missing_value = -9999.f ;
                CV_IMPROAD:vmin = 0.f ;
                CV_IMPROAD:vmax = 0.f ;
                CV_IMPROAD:num_bins = 1 ;
  int NLEV_IMPROAD(numurbl, north_south, east_west) ;
                NLEV_IMPROAD:standard_name = "NLEV_IMPROAD" ;
                NLEV_IMPROAD:units = "" ;
                NLEV_IMPROAD:scale_factor = 1.f ;
                NLEV_IMPROAD:add_offset = 0.f ;
                NLEV_IMPROAD:missing_value = -9999.f ;
                NLEV_IMPROAD:vmin = 0.f ;
                NLEV_IMPROAD:vmax = 0.f ;
                NLEV_IMPROAD:num_bins = 1 ;
  double peatf(north_south, east_west) ;
                peatf:standard_name = "peatf" ;
                peatf:units = "" ;
                peatf:scale_factor = 1.f ;
                peatf:add_offset = 0.f ;
                peatf:missing_value = -9999.f ;
                peatf:vmin = 0.f ;
                peatf:vmax = 0.f ;
                peatf:num_bins = 1 ;
  int abm(north_south, east_west) ;
                abm:standard_name = "abm" ;
                abm:units = "" ;
                abm:scale_factor = 1.f ;
                abm:add_offset = 0.f ;
                abm:missing_value = -9999.f ;
                abm:vmin = 0.f ;
                abm:vmax = 0.f ;
                abm:num_bins = 1 ;
  double gdp(north_south, east_west) ;
                gdp:standard_name = "gdp" ;
                gdp:units = "" ;
                gdp:scale_factor = 1.f ;
                gdp:add_offset = 0.f ;
                gdp:missing_value = -9999.f ;
                gdp:vmin = 0.f ;
                gdp:vmax = 0.f ;
                gdp:num_bins = 1 ;
  double SLOPE(north_south, east_west) ;
                SLOPE:standard_name = "SLOPE" ;
                SLOPE:units = "" ;
                SLOPE:scale_factor = 1.f ;
                SLOPE:add_offset = 0.f ;
                SLOPE:missing_value = -9999.f ;
                SLOPE:vmin = 0.f ;
                SLOPE:vmax = 0.f ;
                SLOPE:num_bins = 1 ;
  double STD_ELEV(north_south, east_west) ;
                STD_ELEV:standard_name = "STD_ELEV" ;
                STD_ELEV:units = "" ;
                STD_ELEV:scale_factor = 1.f ;
                STD_ELEV:add_offset = 0.f ;
                STD_ELEV:missing_value = -9999.f ;
                STD_ELEV:vmin = 0.f ;
                STD_ELEV:vmax = 0.f ;
                STD_ELEV:num_bins = 1 ;
  double binfl(north_south, east_west) ;
                binfl:standard_name = "binfl" ;
                binfl:units = "" ;
                binfl:scale_factor = 1.f ;
                binfl:add_offset = 0.f ;
                binfl:missing_value = -9999.f ;
                binfl:vmin = 0.f ;
                binfl:vmax = 0.f ;
                binfl:num_bins = 1 ;
  double Ws(north_south, east_west) ;
                Ws:standard_name = "Ws" ;
                Ws:units = "" ;
                Ws:scale_factor = 1.f ;
                Ws:add_offset = 0.f ;
                Ws:missing_value = -9999.f ;
                Ws:vmin = 0.f ;
                Ws:vmax = 0.f ;
                Ws:num_bins = 1 ;
  double Dsmax(north_south, east_west) ;
                Dsmax:standard_name = "Dsmax" ;
                Dsmax:units = "" ;
                Dsmax:scale_factor = 1.f ;
                Dsmax:add_offset = 0.f ;
                Dsmax:missing_value = -9999.f ;
                Dsmax:vmin = 0.f ;
                Dsmax:vmax = 0.f ;
                Dsmax:num_bins = 1 ;
  double Ds(north_south, east_west) ;
                Ds:standard_name = "Ds" ;
                Ds:units = "" ;
                Ds:scale_factor = 1.f ;
                Ds:add_offset = 0.f ;
                Ds:missing_value = -9999.f ;
                Ds:vmin = 0.f ;
                Ds:vmax = 0.f ;
                Ds:num_bins = 1 ;
  double LAKEDEPTH(north_south, east_west) ;
                LAKEDEPTH:standard_name = "LAKEDEPTH" ;
                LAKEDEPTH:units = "" ;
                LAKEDEPTH:scale_factor = 1.f ;
                LAKEDEPTH:add_offset = 0.f ;
                LAKEDEPTH:missing_value = -9999.f ;
                LAKEDEPTH:vmin = 0.f ;
                LAKEDEPTH:vmax = 0.f ;
                LAKEDEPTH:num_bins = 1 ;
  double F0(north_south, east_west) ;
                F0:standard_name = "F0" ;
                F0:units = "" ;
                F0:scale_factor = 1.f ;
                F0:add_offset = 0.f ;
                F0:missing_value = -9999.f ;
                F0:vmin = 0.f ;
                F0:vmax = 0.f ;
                F0:num_bins = 1 ;
  double P3(north_south, east_west) ;
                P3:standard_name = "P3" ;
                P3:units = "" ;
                P3:scale_factor = 1.f ;
                P3:add_offset = 0.f ;
                P3:missing_value = -9999.f ;
                P3:vmin = 0.f ;
                P3:vmax = 0.f ;
                P3:num_bins = 1 ;
  double ZWT0(north_south, east_west) ;
                ZWT0:standard_name = "ZWT0" ;
                ZWT0:units = "" ;
                ZWT0:scale_factor = 1.f ;
                ZWT0:add_offset = 0.f ;
                ZWT0:missing_value = -9999.f ;
                ZWT0:vmin = 0.f ;
                ZWT0:vmax = 0.f ;
                ZWT0:num_bins = 1 ;
  double PCT_WETLAND(north_south, east_west) ;
                PCT_WETLAND:standard_name = "PCT_WETLAND" ;
                PCT_WETLAND:units = "" ;
                PCT_WETLAND:scale_factor = 1.f ;
                PCT_WETLAND:add_offset = 0.f ;
                PCT_WETLAND:missing_value = -9999.f ;
                PCT_WETLAND:vmin = 0.f ;
                PCT_WETLAND:vmax = 0.f ;
                PCT_WETLAND:num_bins = 1 ;
  double PCT_LAKE(north_south, east_west) ;
                PCT_LAKE:standard_name = "PCT_LAKE" ;
                PCT_LAKE:units = "" ;
                PCT_LAKE:scale_factor = 1.f ;
                PCT_LAKE:add_offset = 0.f ;
                PCT_LAKE:missing_value = -9999.f ;
                PCT_LAKE:vmin = 0.f ;
                PCT_LAKE:vmax = 0.f ;
                PCT_LAKE:num_bins = 1 ;
  double PCT_GLACIER(north_south, east_west) ;
                PCT_GLACIER:standard_name = "PCT_GLACIER" ;
                PCT_GLACIER:units = "" ;
                PCT_GLACIER:scale_factor = 1.f ;
                PCT_GLACIER:add_offset = 0.f ;
                PCT_GLACIER:missing_value = -9999.f ;
                PCT_GLACIER:vmin = 0.f ;
                PCT_GLACIER:vmax = 0.f ;
                PCT_GLACIER:num_bins = 1 ;
  double GLC_MEC(nglcecp1) ;
                GLC_MEC:standard_name = "GLC_MEC" ;
                GLC_MEC:units = "" ;
                GLC_MEC:scale_factor = 1.f ;
                GLC_MEC:add_offset = 0.f ;
                GLC_MEC:missing_value = -9999.f ;
                GLC_MEC:vmin = 0.f ;
                GLC_MEC:vmax = 0.f ;
                GLC_MEC:num_bins = 1 ;
  double PCT_GLC_MEC(nglcec, north_south, east_west) ;
                PCT_GLC_MEC:standard_name = "PCT_GLC_MEC" ;
                PCT_GLC_MEC:units = "" ;
                PCT_GLC_MEC:scale_factor = 1.f ;
                PCT_GLC_MEC:add_offset = 0.f ;
                PCT_GLC_MEC:missing_value = -9999.f ;
                PCT_GLC_MEC:vmin = 0.f ;
                PCT_GLC_MEC:vmax = 0.f ;
                PCT_GLC_MEC:num_bins = 1 ;
  double PCT_GLC_MEC_GIC(nglcec, north_south, east_west) ;
                PCT_GLC_MEC_GIC:standard_name = "PCT_GLC_MEC_GIC" ;
                PCT_GLC_MEC_GIC:units = "" ;
                PCT_GLC_MEC_GIC:scale_factor = 1.f ;
                PCT_GLC_MEC_GIC:add_offset = 0.f ;
                PCT_GLC_MEC_GIC:missing_value = -9999.f ;
                PCT_GLC_MEC_GIC:vmin = 0.f ;
                PCT_GLC_MEC_GIC:vmax = 0.f ;
                PCT_GLC_MEC_GIC:num_bins = 1 ;
  double PCT_GLC_MEC_ICESHEET(nglcec, north_south, east_west) ;
                PCT_GLC_MEC_ICESHEET:standard_name = "PCT_GLC_MEC_ICESHEET" ;
                PCT_GLC_MEC_ICESHEET:units = "" ;
                PCT_GLC_MEC_ICESHEET:scale_factor = 1.f ;
                PCT_GLC_MEC_ICESHEET:add_offset = 0.f ;
                PCT_GLC_MEC_ICESHEET:missing_value = -9999.f ;
                PCT_GLC_MEC_ICESHEET:vmin = 0.f ;
                PCT_GLC_MEC_ICESHEET:vmax = 0.f ;
                PCT_GLC_MEC_ICESHEET:num_bins = 1 ;
  double PCT_GLC_GIC(north_south, east_west) ;
                PCT_GLC_GIC:standard_name = "PCT_GLC_GIC" ;
                PCT_GLC_GIC:units = "" ;
                PCT_GLC_GIC:scale_factor = 1.f ;
                PCT_GLC_GIC:add_offset = 0.f ;
                PCT_GLC_GIC:missing_value = -9999.f ;
                PCT_GLC_GIC:vmin = 0.f ;
                PCT_GLC_GIC:vmax = 0.f ;
                PCT_GLC_GIC:num_bins = 1 ;
  double PCT_GLC_ICESHEET(north_south, east_west) ;
                PCT_GLC_ICESHEET:standard_name = "PCT_GLC_ICESHEET" ;
                PCT_GLC_ICESHEET:units = "" ;
                PCT_GLC_ICESHEET:scale_factor = 1.f ;
                PCT_GLC_ICESHEET:add_offset = 0.f ;
                PCT_GLC_ICESHEET:missing_value = -9999.f ;
                PCT_GLC_ICESHEET:vmin = 0.f ;
                PCT_GLC_ICESHEET:vmax = 0.f ;
                PCT_GLC_ICESHEET:num_bins = 1 ;
  double TOPO_GLC_MEC(nglcec, north_south, east_west) ;
                TOPO_GLC_MEC:standard_name = "TOPO_GLC_MEC" ;
                TOPO_GLC_MEC:units = "" ;
                TOPO_GLC_MEC:scale_factor = 1.f ;
                TOPO_GLC_MEC:add_offset = 0.f ;
                TOPO_GLC_MEC:missing_value = -9999.f ;
                TOPO_GLC_MEC:vmin = 0.f ;
                TOPO_GLC_MEC:vmax = 0.f ;
                TOPO_GLC_MEC:num_bins = 1 ;
  double TOPO(north_south, east_west) ;
                TOPO:standard_name = "TOPO" ;
                TOPO:units = "" ;
                TOPO:scale_factor = 1.f ;
                TOPO:add_offset = 0.f ;
                TOPO:missing_value = -9999.f ;
                TOPO:vmin = 0.f ;
                TOPO:vmax = 0.f ;
                TOPO:num_bins = 1 ;
  double PCT_URBAN(numurbl, north_south, east_west) ;
                PCT_URBAN:standard_name = "PCT_URBAN" ;
                PCT_URBAN:units = "" ;
                PCT_URBAN:scale_factor = 1.f ;
                PCT_URBAN:add_offset = 0.f ;
                PCT_URBAN:missing_value = -9999.f ;
                PCT_URBAN:vmin = 0.f ;
                PCT_URBAN:vmax = 0.f ;
                PCT_URBAN:num_bins = 1 ;
  int URBAN_REGION_ID(north_south, east_west) ;
                URBAN_REGION_ID:standard_name = "URBAN_REGION_ID" ;
                URBAN_REGION_ID:units = "" ;
                URBAN_REGION_ID:scale_factor = 1.f ;
                URBAN_REGION_ID:add_offset = 0.f ;
                URBAN_REGION_ID:missing_value = -9999.f ;
                URBAN_REGION_ID:vmin = 0.f ;
                URBAN_REGION_ID:vmax = 0.f ;
                URBAN_REGION_ID:num_bins = 1 ;
// global attributes:
		:MAP_PROJECTION = "EQUIDISTANT CYLINDRICAL" ;
		:SOUTH_WEST_CORNER_LAT = -90.0f ;
		:SOUTH_WEST_CORNER_LON = 0.0f ;
		:DX = 1.25f ;
		:DY = 0.942f ;
		:INC_WATER_PTS = "false" ;
		:LANDCOVER_SCHEME = "UMD" ;
		:BARESOILCLASS = 12 ;
		:URBANCLASS = 13 ;
		:SNOWCLASS = 0 ;
		:WATERCLASS = 14 ;
		:WETLANDCLASS = 0 ;
		:GLACIERCLASS = 0 ;
		:NUMVEGTYPES = 13 ;
		:LANDMASK_SOURCE = "AVHRR" ;
		:SFCMODELS = "CLM.4.5" ;
		:SOILTEXT_SCHEME = "Soil texture not selected" ;
		:LAISAI_DATA_INTERVAL = "monthly" ;
		:title = "Land Data Toolkit (LDT) parameter-processed output" ;
		:institution = "NASA GSFC Hydrological Sciences Laboratory" ;
		:history = "created on date: 2015-09-14T12:32:09.195" ;
		:references = "Kumar_etal_EMS_2006, Peters-Lidard_etal_ISSE_2007" ;
		:comment = "website: http://lis.gsfc.nasa.gov/" ;
